module qe(i, q, y15,y14,y13,y12,y11,y10,y9,y8,y7,y6,y5,y4,y3,y2,y1);
   input i, q;

   output y15,y14,y13,y12,y11,y10,y9,y8,y7,y6,y5,y4,y3,y2,y1;

   


endmodule
