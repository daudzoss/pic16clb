module terminator(y0,y1,y2,y3);
input y3,y2,y1,y0;
wire w3,w2,w1,w0;
assign w3 = y3;
assign w2 = y2;
assign w1 = y1;
assign w0 = y0;
endmodule